`include "uvm_macros.svh"
import uvm_pkg::*;
`include "seq_item.sv"
`include "sequence.sv"
`include "callback.sv"
`include "master_sequencer.sv"
`include "slave_sequencer.sv"
`include "interface.sv"
`include "master_driver.sv"
`include "slave_driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "top.sv"
